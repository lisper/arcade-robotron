library IEEE;
   use IEEE.std_logic_1164.all;
   use IEEE.std_logic_arith.all;
library unisim;
   use unisim.vcomponents.all;
   
entity ROM_SND_F000 is
   port(
      clk    : in  std_logic;
      rst    : in  std_logic;
      cs     : in  std_logic;
      addr   : in  std_logic_vector(10 downto 0);
      data   : out std_logic_vector(7 downto 0)
   );
end ROM_SND_F000;

architecture rtl of ROM_SND_F000 is
   signal dp : std_logic;
begin
   ROM: RAMB16_S9
      generic map (
         INIT_00 => x"008e0f5343494e4f525443454c4520534d41494c4c4957203238393129432876",
         INIT_01 => x"970197009703974f059701a73c8603a73786026f00a7ff86036f016f0004ce7f",
         INIT_02 => x"271a007afd265a5c54545406d6092a15d6808607dfebf0ce0cdffe200e049702",
         INIT_03 => x"d70bcb06db5806d61dd77fc4db2715d6df261d007a4c271c007a4c271b007a4c",
         INIT_04 => x"19d405207fc419d4062b06d607df4e27e4f08c0907de2dd721d60e262d007a06",
         INIT_05 => x"186a1227186d1400ce03201300ce08201200cea22000ad07de32161b36507fc4",
         INIT_06 => x"4ff07e00ad07de16046004ab08e700e600e7122714e110eb00e618e70ce60e26",
         INIT_07 => x"f220eef3ce3946f0bd65f9bd1cc6d2f3ce390004f75454545454545454390cde",
         INIT_08 => x"028000a66000ced92096f4cede207af4cee32042f4cee82026f4ceed200af4ce",
         INIT_09 => x"000473fd260912df0812de00047f14df8003ce12df0100ce49f37e30f3bd00a7",
         INIT_0a => x"17df16974400ce0186058de0ffce208614dfc0fece1297ff86eb20fd260914de",
         INIT_0b => x"de14007c03241597169b1596ef26091297149912961397159b1396218d1000ce",
         INIT_0c => x"fd264a028612d6f92420800004b7e086098df924208b0004b74f39db26179c14",
         INIT_0d => x"d88b44444419971c9b1996fd264a1286109780861a97f1861c97808639f8265a",
         INIT_0e => x"d0c6bcb0a5988c8039d52620811c961c007ae22610007a0004b700a61ade1b97",
         INIT_0f => x"2f39434f5a6773808c98a5b0bcc6d0dae2eaf0f5fafdfefffefdfaf5f0eae2da",
         INIT_10 => x"14df5ff2ce02047f73675a4f43392f251d150f0a050201000102050a0f151d25",
         INIT_11 => x"0500ce12960004b713960fc4129714df080801e613d7f0c401e6332700a614de",
         INIT_12 => x"01390204b78086c720df265af7264afd26090500ce129600047ff7264afd2609",
         INIT_13 => x"2e007a0000f1c0f1a0f180f160f140f220f410f40cf408f806f804f803fc02fc",
         INIT_14 => x"12007a1727090004b71200f7202709c001ce2ed69f86139704862ed7a0c60420",
         INIT_15 => x"862ed711c639d42210c113d0dd20f82612007a07270900047312d70f2709f826",
         INIT_16 => x"ceeb8dbef4ce09d7ffc6f420b8f4ce3949f3bd30f3bd2620b2f4cec5201397fe",
         INIT_17 => x"86f120dcf4ce0997ff86fa20308dd88dd6f4cedd20caf4ce39f3265ae68dc4f4",
         INIT_18 => x"298d13970c8b444406970b8b069b480696218de2f4ce30c6e820d0f4ce0997ff",
         INIT_19 => x"169703a6159702a6149701a6139700a6393232390997032a0880099639ec265a",
         INIT_1a => x"13d643fd265a0004b713d6431ad714d619d717d637099639189705a6179704a6",
         INIT_1b => x"13d619d70004b717d643de2619007a16271a007afd265a0004b7090809080020",
         INIT_1c => x"05c013d7062716d116d115d013d61ad70004b714d6430109081520011e2b189b",
         INIT_1d => x"171a1c2520272c3346503e3a00f9f6f900070a078026012680daffda3933b820",
         INIT_1e => x"ffff90ffffffffffffff90ffffff0070321e0a06050403020102030833101114",
         INIT_1f => x"0181000008010000014800003f3f000001480000000000000000ffffffffffff",
         INIT_20 => x"ff3100000101000005050000100100003f3f00001001000008010000ff010000",
         INIT_21 => x"0001000000020000007f00000001000000300000007f00000030000005050000",
         INIT_22 => x"680ca00000ff0000000000000000a00000ff040000047f00007f040000040000",
         INIT_23 => x"7f3f0000040100ffffff000000000000000000ffffff0080800c000f1f070068",
         INIT_24 => x"80027f007f0a300080020000ff0500000048000000010000ff05000004010000",
         INIT_25 => x"032000ff80ff030100ffc30201ff000080c0000010c015001001200080c03000",
         INIT_26 => x"100201e000ff0c01024800ff0c01034800ff040204fe00ff2001035000ff50ff",
         INIT_27 => x"09c692fbbd08fcce0edf1200ce1b4848481600ff060102ff80600000ff5000ff",
         INIT_28 => x"000473fa264a1027090004731b9617de1c9713961b9712960004b71a9665f97e",
         INIT_29 => x"97159b1c961b97149b1b960004b7008b43012b0004b6e820fa264a0527091c96",
         INIT_2a => x"03c6199701861220ffc660861997ff8639b9261297129b06271996cb2616911c",
         INIT_2b => x"76440698444444069614d614d70004b7ff861897002010c6c0861997fe860a20",
         INIT_2c => x"971497208639db261897199b1896e5265afd264a189600047303240600760500",
         INIT_2d => x"060076050076440698444444069614d613d715df12970020ffc60100ce018617",
         INIT_2e => x"cc20d02717960815de092712d013d6e1265afd260915de0004b7139602240086",
         INIT_2f => x"dbf67e33f6bd2ef6cecef6bd33f6bd29f6ce05df00a5ce2af7bd23df00f6ce39",
         INIT_30 => x"20ac58140230c02820ff54e954080220ee60100232d03014ff40b44014021090",
         INIT_31 => x"a6129702a6139701a62a9700a6010001fc300100fc1030002218ff58a6580802",
         INIT_32 => x"007d5c8d388d2d8d0004f759f8262f912e96588d308de98d392f9704a6179703",
         INIT_33 => x"9614007fd0202e007a2f007ad8202f007c052bdf2717007de42614007de42713",
         INIT_34 => x"24008606007605007644289639078408289706984444440696392d007f2e972f",
         INIT_35 => x"042714912a963914007c542dd62e970820090804272e007a2f96392d97139602",
         INIT_36 => x"bda88d9f8d27007f22970e862b007f21007f3913971290139614007f09200908",
         INIT_37 => x"22007a2696e220528d6d8d1d8d718d0a8d758dcd8d798dbd8d64f7bdb08d64f7",
         INIT_38 => x"7f29202a261396080727299121963921972b9b2196229768200a261300b60727",
         INIT_39 => x"299704a6269703a62c9702a6259701a61727209700a623de27007f2b007f2100",
         INIT_3a => x"962197259620007f390908032004261391062720963932323923df92fbbd0586",
         INIT_3b => x"25208bf7ce2a2085f7ce00d701c6390004b71b43012a2797219b2796392b972c",
         INIT_3c => x"018001001040010101e803ff010001000003000000000001000000202091f7ce",
         INIT_3d => x"04b616de14007f16df12d7189704ee03e602a6159701a6199700a697f7ceff40",
         INIT_3e => x"22069114d613d715db05d4042719007d12d60600760500765406d85454541600",
         INIT_3f => x"910425139214d00004b71427091020f02306911625139914db0004b726270912"
      )
      port map (
         do    => data,
         dop(0)  => dp,
         addr    => addr,
         clk     => clk,
         di      => "00000000",
         dip(0)  => '0',
         en      => cs,
         ssr     => rst,
         we      => '0'
      );
end architecture rtl;

library IEEE;
   use IEEE.std_logic_1164.all;
   use IEEE.std_logic_arith.all;
library unisim;
   use unisim.vcomponents.all;
   
entity ROM_SND_F800 is
   port(
      clk    : in  std_logic;
      rst    : in  std_logic;
      cs     : in  std_logic;
      addr   : in  std_logic_vector(10 downto 0);
      data   : out std_logic_vector(7 downto 0)
   );
end ROM_SND_F800;

architecture rtl of ROM_SND_F800 is
   signal dp : std_logic;
begin
   ROM: RAMB16_S9
      generic map (
         INIT_00 => x"129914dbff82504356445644564414d61296b32718d6b7200004b70696f02206",
         INIT_01 => x"04250ade10970a9910960bdb0adf6400ce0e97fc8639922607c19626129714d7",
         INIT_02 => x"4f10970004b74f39dc200004b700a60ede0f97478b0f840adf11270803200020",
         INIT_03 => x"008c08006f1200ce39e82a10007c000473f12a4cfd265a12c600047303261091",
         INIT_04 => x"008c080810007410db022a01a700ab01a65f109780861200ce12974086f8261a",
         INIT_05 => x"08085c006a02e741c6042637810b2700a65f1200cedc2611007c0004f7ec261a",
         INIT_06 => x"007a2d2700a657fcce109704007f7ffb7e038d3904007a39bf265dea261a008c",
         INIT_07 => x"de0e8d12df02ee01a6149700a60ede0cdf92fbbd0edf08f12092fbbd4c062710",
         INIT_08 => x"2002800800e701c609270381152302801500ce3939e8260c9c0edf080808080e",
         INIT_09 => x"14d411d75c1100f64f12de02e737c601e7f9c600e77ec60808016f00e791c6f1",
         INIT_0a => x"27090004b748484848481b008954008954008954008954008954008954008954",
         INIT_0b => x"7f39019700974f3932ef265a080cde0edf0800a70ede0cdf00a6363915007e03",
         INIT_0c => x"bd16007c94fabd4348480196dcf9bd0e863901974c4f01261d817f8401960000",
         INIT_0d => x"f7204a0ecb052314815f10208602d75c5f01261fc102d6eef4bd0386f82096fa",
         INIT_0e => x"1b1b581689fa7e6920058d0d8603007c09260396fb2003f5bd12d7fb264a05cb",
         INIT_0f => x"970f8414d7545454541601a612d75454545413970f841600a692fbbd45fece1b",
         INIT_10 => x"fabd199702a60aded0fabd17dff32092fbbd4c00a6082b10007a32fdce0adf10",
         INIT_11 => x"df92fbbd22007f1adf1792fbbd02ffce06a61605a6169704a6159703a60adee2",
         INIT_12 => x"20962300ce0cdf0813d626271c9c2097229b00a60cde0cdf1ade21971296391c",
         INIT_13 => x"628d1496df2001010908090809080908da275af1261e9c080004b700a6fd264a",
         INIT_14 => x"062b15007d22965f1ade2297229b3d2716007a4227159646260396c12621007a",
         INIT_15 => x"3901265ddd261c9c085c1adf03265d0f2008275d0525022700ab0b20082500ab",
         INIT_16 => x"df0ede65f9bd0800e617de0edf2300ce3942fa7e168d1996088d062714961cdf",
         INIT_17 => x"de0cdf085454545401e610d711d60cde0edf11972300ce0cdf17de2b274d391e",
         INIT_18 => x"df1200ce07dfebf0ce0204b67f008e39de261e9c0800a7fa2610007a1000a60e",
         INIT_19 => x"3f274d03d70227128102d702270e815fcdf8bd032704d63f84430e09d7afc60e",
         INIT_1a => x"dcf9bd08220c8112201c80242039800c20108008222a81082e3d81142d1f814a",
         INIT_1b => x"9603f5bdeef4bd1c80082000ad00ee218dc4fbce480d800e221b811a2042fabd",
         INIT_1c => x"390cde0c007c03240d970d9b0cdf8ff97e72f77e0327009603974ffe27019a00",
         INIT_1d => x"bd0186d2f8bd0286a2f7bd3e012700e1f82600f08c0900e95fffffce7f008e0f",
         INIT_1e => x"c9f878f859f82bf880f77bf762f59bf579f9ccf95af57ff972f7a4f9dc20d2f8",
         INIT_1f => x"e1f550f514f10ff128f1bbf208f3fff2e8f2d6f2d1f2f6f2eff00af1fbf00cf9",
         INIT_20 => x"0201fc008128ffff00028108000128ffff8000e110000140a2f7a4f147f118f2",
         INIT_21 => x"0160fffc000201fc008128ff00800468ff08ff00ff00800441180001fffffc00",
         INIT_22 => x"55050400550504f81c8c5bb640bf49a47373a449bf40b65b8c80fe0002e10857",
         INIT_23 => x"041d3e66060400cb041d1fb0413b17f855050400550504f855050400550504f8",
         INIT_24 => x"041df866060400cb041d7cfe1f040097033f7c6606040097033f3efe1f0400cb",
         INIT_25 => x"05127ccb041d7c97033f7cca2c040097033ff86606040097033f7c66060400cb",
         INIT_26 => x"03373ecb041d7c6105127cb3050d7c6606047cb3050d7c6105127cb3050d7c61",
         INIT_27 => x"05127ccb041d7c8604237ccb041d7c6105127cb3050d7c6606047c97033f3ece",
         INIT_28 => x"1f040097033f7c6606040097033f3e66060400cb041d7c66060400cb041d3e61",
         INIT_29 => x"00804000082400247fd9ffd97f0804080d12171d232930373f4700ee2f1df8fe",
         INIT_2a => x"947f6a6d8dbfe7ecc57f104e24090009244e7fb0d9f5fff5d9b07f10408000ff",
         INIT_2b => x"d1c8bfb5aba0958a4800000000ffffffff00000000ffffffff10391217407192",
         INIT_2c => x"545f6a757f8a95a0abb5bfc8d1dae1e8eef3f7fbfdfefffefdfbf7f3eee8e1da",
         INIT_2d => x"7f756a5f544a40372e251e17110c0804020100010204080c11171e252e37404a",
         INIT_2e => x"9dd0b8ff761000000000ffffffff0837190600061937597b98acb3ac987b5910",
         INIT_2f => x"504b45480000f400e800dc00e200dc00e800f4001063329c4e8681ea76826ae6",
         INIT_30 => x"454b50565b6064696d7174777a7c7e7f7f807f7f7e7c7a7774716d6964605b56",
         INIT_31 => x"25201c17130f0c090604020101000101020406090c0f13171c20252a30353b40",
         INIT_32 => x"0d000100311147010f011105116d2700ff1a051231160000002481403b35302a",
         INIT_33 => x"001131690100fd0000151b0d00ff1135215b0f0000004541471400000012f41b",
         INIT_34 => x"690410ff00121f9a06020002106a940602000353f6470101010115016a030001",
         INIT_35 => x"010030210d0e00000011f40d0e0000001714280901ff000612000d00ff001131",
         INIT_36 => x"21df1600000019f2c6180000002282b31200000018f4a40900ff0010131b0d00",
         INIT_37 => x"00ff1115036d270000d002416a030001001931a40e00000019f10d1b00ff0030",
         INIT_38 => x"020101e0c0603010100808040402020101404450586068707880889098a01b0d",
         INIT_39 => x"38302820100808040402020101807c78747074787c800c0a0908070605040302",
         INIT_3a => x"0402014008400840084008400840084008400840084008c0b0a0807060504840",
         INIT_3b => x"14100c0a0806050404030302020101010101081040161412100f0e0c0b0a0908",
         INIT_3c => x"1a191817080c0a09080701010102020304050607080a0c102030405040302018",
         INIT_3d => x"0801100801100801100801004840503058286020701878108008000000001c1b",
         INIT_3e => x"4020104020104020104020104020104020104020104020100010080110080110",
         INIT_3f => x"1df0a0fb1df011fb004b0b4a0a49094808470746064505440443034202400100"
      )
      port map (
         do    => data,
         dop(0)  => dp,
         addr    => addr,
         clk     => clk,
         di      => "00000000",
         dip(0)  => '0',
         en      => cs,
         ssr     => rst,
         we      => '0'
      );
end architecture rtl;

